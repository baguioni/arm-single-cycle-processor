module plus_4(input [31:0] number, output [31:0] number_plus_4);
	assign number_plus_4 = number + 4;
endmodule
